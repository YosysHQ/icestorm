module top (input C, D, output Q);
	SB_DFF ff (.C(C), .D(D), .Q(Q));
endmodule
